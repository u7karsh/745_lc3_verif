// Data memory
typedef reg[15:0] data_t;

typedef enum {
   WARN,
   FATAL
} severityT;
